library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity nbitregbank is
    generic (n: natural:=8);
    port(
        wr_data_reg: in std_lo
    )